/RAID2/COURSE/iclab/iclabTA01/UMC018_CBDK/CIC/SOCE/lef/BONDPAD.lef