../02_SYN/Netlist/Program_Wrapper.sv