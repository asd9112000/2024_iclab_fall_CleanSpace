/RAID2/COURSE/iclab/iclabTA01/UMC018_CBDK/CIC/SOCE/lef/fsa0m_a_generic_core.lef