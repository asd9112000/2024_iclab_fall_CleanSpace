/RAID2/COURSE/iclab/iclabTA05/TA_Lab09/Exercise/01_RTL/Program.sv