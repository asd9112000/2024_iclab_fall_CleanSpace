/RAID2/COURSE/BackUp/2023_Spring/iclab/iclabta01/LAB10_TA_DESIGN_24A/TA_Program.sv