/RAID2/COURSE/iclab/iclabTA01/UMC018_CBDK/CIC/SOCE/lef/header6_V55_20ka_cic.lef