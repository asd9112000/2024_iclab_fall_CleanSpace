# 
#              Synchronous Dual Port SRAM Compiler 
# 
#                    UMC 0.18um Generic Logic Process 
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : W1024_B8_BM2
#       Words            : 1024
#       Bits             : 8
#       Byte-Write       : 1
#       Aspect Ratio     : 2
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2024/10/07 09:38:09
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO W1024_B8_BM2
CLASS BLOCK ;
FOREIGN W1024_B8_BM2 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 544.980 BY 350.000 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME5 ;
  RECT 543.860 336.900 544.980 340.140 ;
  LAYER ME4 ;
  RECT 543.860 336.900 544.980 340.140 ;
  LAYER ME3 ;
  RECT 543.860 336.900 544.980 340.140 ;
  LAYER ME2 ;
  RECT 543.860 336.900 544.980 340.140 ;
  LAYER ME1 ;
  RECT 543.860 336.900 544.980 340.140 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 329.060 544.980 332.300 ;
  LAYER ME4 ;
  RECT 543.860 329.060 544.980 332.300 ;
  LAYER ME3 ;
  RECT 543.860 329.060 544.980 332.300 ;
  LAYER ME2 ;
  RECT 543.860 329.060 544.980 332.300 ;
  LAYER ME1 ;
  RECT 543.860 329.060 544.980 332.300 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 321.220 544.980 324.460 ;
  LAYER ME4 ;
  RECT 543.860 321.220 544.980 324.460 ;
  LAYER ME3 ;
  RECT 543.860 321.220 544.980 324.460 ;
  LAYER ME2 ;
  RECT 543.860 321.220 544.980 324.460 ;
  LAYER ME1 ;
  RECT 543.860 321.220 544.980 324.460 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 282.020 544.980 285.260 ;
  LAYER ME4 ;
  RECT 543.860 282.020 544.980 285.260 ;
  LAYER ME3 ;
  RECT 543.860 282.020 544.980 285.260 ;
  LAYER ME2 ;
  RECT 543.860 282.020 544.980 285.260 ;
  LAYER ME1 ;
  RECT 543.860 282.020 544.980 285.260 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 274.180 544.980 277.420 ;
  LAYER ME4 ;
  RECT 543.860 274.180 544.980 277.420 ;
  LAYER ME3 ;
  RECT 543.860 274.180 544.980 277.420 ;
  LAYER ME2 ;
  RECT 543.860 274.180 544.980 277.420 ;
  LAYER ME1 ;
  RECT 543.860 274.180 544.980 277.420 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 266.340 544.980 269.580 ;
  LAYER ME4 ;
  RECT 543.860 266.340 544.980 269.580 ;
  LAYER ME3 ;
  RECT 543.860 266.340 544.980 269.580 ;
  LAYER ME2 ;
  RECT 543.860 266.340 544.980 269.580 ;
  LAYER ME1 ;
  RECT 543.860 266.340 544.980 269.580 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 258.500 544.980 261.740 ;
  LAYER ME4 ;
  RECT 543.860 258.500 544.980 261.740 ;
  LAYER ME3 ;
  RECT 543.860 258.500 544.980 261.740 ;
  LAYER ME2 ;
  RECT 543.860 258.500 544.980 261.740 ;
  LAYER ME1 ;
  RECT 543.860 258.500 544.980 261.740 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 250.660 544.980 253.900 ;
  LAYER ME4 ;
  RECT 543.860 250.660 544.980 253.900 ;
  LAYER ME3 ;
  RECT 543.860 250.660 544.980 253.900 ;
  LAYER ME2 ;
  RECT 543.860 250.660 544.980 253.900 ;
  LAYER ME1 ;
  RECT 543.860 250.660 544.980 253.900 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 242.820 544.980 246.060 ;
  LAYER ME4 ;
  RECT 543.860 242.820 544.980 246.060 ;
  LAYER ME3 ;
  RECT 543.860 242.820 544.980 246.060 ;
  LAYER ME2 ;
  RECT 543.860 242.820 544.980 246.060 ;
  LAYER ME1 ;
  RECT 543.860 242.820 544.980 246.060 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 203.620 544.980 206.860 ;
  LAYER ME4 ;
  RECT 543.860 203.620 544.980 206.860 ;
  LAYER ME3 ;
  RECT 543.860 203.620 544.980 206.860 ;
  LAYER ME2 ;
  RECT 543.860 203.620 544.980 206.860 ;
  LAYER ME1 ;
  RECT 543.860 203.620 544.980 206.860 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 195.780 544.980 199.020 ;
  LAYER ME4 ;
  RECT 543.860 195.780 544.980 199.020 ;
  LAYER ME3 ;
  RECT 543.860 195.780 544.980 199.020 ;
  LAYER ME2 ;
  RECT 543.860 195.780 544.980 199.020 ;
  LAYER ME1 ;
  RECT 543.860 195.780 544.980 199.020 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 187.940 544.980 191.180 ;
  LAYER ME4 ;
  RECT 543.860 187.940 544.980 191.180 ;
  LAYER ME3 ;
  RECT 543.860 187.940 544.980 191.180 ;
  LAYER ME2 ;
  RECT 543.860 187.940 544.980 191.180 ;
  LAYER ME1 ;
  RECT 543.860 187.940 544.980 191.180 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 180.100 544.980 183.340 ;
  LAYER ME4 ;
  RECT 543.860 180.100 544.980 183.340 ;
  LAYER ME3 ;
  RECT 543.860 180.100 544.980 183.340 ;
  LAYER ME2 ;
  RECT 543.860 180.100 544.980 183.340 ;
  LAYER ME1 ;
  RECT 543.860 180.100 544.980 183.340 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 172.260 544.980 175.500 ;
  LAYER ME4 ;
  RECT 543.860 172.260 544.980 175.500 ;
  LAYER ME3 ;
  RECT 543.860 172.260 544.980 175.500 ;
  LAYER ME2 ;
  RECT 543.860 172.260 544.980 175.500 ;
  LAYER ME1 ;
  RECT 543.860 172.260 544.980 175.500 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 164.420 544.980 167.660 ;
  LAYER ME4 ;
  RECT 543.860 164.420 544.980 167.660 ;
  LAYER ME3 ;
  RECT 543.860 164.420 544.980 167.660 ;
  LAYER ME2 ;
  RECT 543.860 164.420 544.980 167.660 ;
  LAYER ME1 ;
  RECT 543.860 164.420 544.980 167.660 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 125.220 544.980 128.460 ;
  LAYER ME4 ;
  RECT 543.860 125.220 544.980 128.460 ;
  LAYER ME3 ;
  RECT 543.860 125.220 544.980 128.460 ;
  LAYER ME2 ;
  RECT 543.860 125.220 544.980 128.460 ;
  LAYER ME1 ;
  RECT 543.860 125.220 544.980 128.460 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 117.380 544.980 120.620 ;
  LAYER ME4 ;
  RECT 543.860 117.380 544.980 120.620 ;
  LAYER ME3 ;
  RECT 543.860 117.380 544.980 120.620 ;
  LAYER ME2 ;
  RECT 543.860 117.380 544.980 120.620 ;
  LAYER ME1 ;
  RECT 543.860 117.380 544.980 120.620 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 109.540 544.980 112.780 ;
  LAYER ME4 ;
  RECT 543.860 109.540 544.980 112.780 ;
  LAYER ME3 ;
  RECT 543.860 109.540 544.980 112.780 ;
  LAYER ME2 ;
  RECT 543.860 109.540 544.980 112.780 ;
  LAYER ME1 ;
  RECT 543.860 109.540 544.980 112.780 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 101.700 544.980 104.940 ;
  LAYER ME4 ;
  RECT 543.860 101.700 544.980 104.940 ;
  LAYER ME3 ;
  RECT 543.860 101.700 544.980 104.940 ;
  LAYER ME2 ;
  RECT 543.860 101.700 544.980 104.940 ;
  LAYER ME1 ;
  RECT 543.860 101.700 544.980 104.940 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 93.860 544.980 97.100 ;
  LAYER ME4 ;
  RECT 543.860 93.860 544.980 97.100 ;
  LAYER ME3 ;
  RECT 543.860 93.860 544.980 97.100 ;
  LAYER ME2 ;
  RECT 543.860 93.860 544.980 97.100 ;
  LAYER ME1 ;
  RECT 543.860 93.860 544.980 97.100 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 86.020 544.980 89.260 ;
  LAYER ME4 ;
  RECT 543.860 86.020 544.980 89.260 ;
  LAYER ME3 ;
  RECT 543.860 86.020 544.980 89.260 ;
  LAYER ME2 ;
  RECT 543.860 86.020 544.980 89.260 ;
  LAYER ME1 ;
  RECT 543.860 86.020 544.980 89.260 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 46.820 544.980 50.060 ;
  LAYER ME4 ;
  RECT 543.860 46.820 544.980 50.060 ;
  LAYER ME3 ;
  RECT 543.860 46.820 544.980 50.060 ;
  LAYER ME2 ;
  RECT 543.860 46.820 544.980 50.060 ;
  LAYER ME1 ;
  RECT 543.860 46.820 544.980 50.060 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 38.980 544.980 42.220 ;
  LAYER ME4 ;
  RECT 543.860 38.980 544.980 42.220 ;
  LAYER ME3 ;
  RECT 543.860 38.980 544.980 42.220 ;
  LAYER ME2 ;
  RECT 543.860 38.980 544.980 42.220 ;
  LAYER ME1 ;
  RECT 543.860 38.980 544.980 42.220 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 31.140 544.980 34.380 ;
  LAYER ME4 ;
  RECT 543.860 31.140 544.980 34.380 ;
  LAYER ME3 ;
  RECT 543.860 31.140 544.980 34.380 ;
  LAYER ME2 ;
  RECT 543.860 31.140 544.980 34.380 ;
  LAYER ME1 ;
  RECT 543.860 31.140 544.980 34.380 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 23.300 544.980 26.540 ;
  LAYER ME4 ;
  RECT 543.860 23.300 544.980 26.540 ;
  LAYER ME3 ;
  RECT 543.860 23.300 544.980 26.540 ;
  LAYER ME2 ;
  RECT 543.860 23.300 544.980 26.540 ;
  LAYER ME1 ;
  RECT 543.860 23.300 544.980 26.540 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 15.460 544.980 18.700 ;
  LAYER ME4 ;
  RECT 543.860 15.460 544.980 18.700 ;
  LAYER ME3 ;
  RECT 543.860 15.460 544.980 18.700 ;
  LAYER ME2 ;
  RECT 543.860 15.460 544.980 18.700 ;
  LAYER ME1 ;
  RECT 543.860 15.460 544.980 18.700 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 7.620 544.980 10.860 ;
  LAYER ME4 ;
  RECT 543.860 7.620 544.980 10.860 ;
  LAYER ME3 ;
  RECT 543.860 7.620 544.980 10.860 ;
  LAYER ME2 ;
  RECT 543.860 7.620 544.980 10.860 ;
  LAYER ME1 ;
  RECT 543.860 7.620 544.980 10.860 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER ME4 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER ME3 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER ME2 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER ME1 ;
  RECT 0.000 336.900 1.120 340.140 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER ME4 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER ME3 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER ME2 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER ME1 ;
  RECT 0.000 329.060 1.120 332.300 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER ME4 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER ME3 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER ME2 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER ME1 ;
  RECT 0.000 321.220 1.120 324.460 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER ME4 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER ME3 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER ME2 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER ME1 ;
  RECT 0.000 282.020 1.120 285.260 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER ME4 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER ME3 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER ME2 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER ME1 ;
  RECT 0.000 274.180 1.120 277.420 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER ME4 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER ME3 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER ME2 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER ME1 ;
  RECT 0.000 266.340 1.120 269.580 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER ME4 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER ME3 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER ME2 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER ME1 ;
  RECT 0.000 258.500 1.120 261.740 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER ME4 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER ME3 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER ME2 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER ME1 ;
  RECT 0.000 250.660 1.120 253.900 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER ME4 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER ME3 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER ME2 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER ME1 ;
  RECT 0.000 242.820 1.120 246.060 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER ME4 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER ME3 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER ME2 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER ME1 ;
  RECT 0.000 203.620 1.120 206.860 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER ME4 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER ME3 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER ME2 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER ME1 ;
  RECT 0.000 195.780 1.120 199.020 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER ME4 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER ME3 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER ME2 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER ME1 ;
  RECT 0.000 187.940 1.120 191.180 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER ME4 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER ME3 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER ME2 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER ME1 ;
  RECT 0.000 180.100 1.120 183.340 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER ME4 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER ME3 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER ME2 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER ME1 ;
  RECT 0.000 172.260 1.120 175.500 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER ME4 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER ME3 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER ME2 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER ME1 ;
  RECT 0.000 164.420 1.120 167.660 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER ME4 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER ME3 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER ME2 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER ME1 ;
  RECT 0.000 125.220 1.120 128.460 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER ME4 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER ME3 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER ME2 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER ME1 ;
  RECT 0.000 117.380 1.120 120.620 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER ME4 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER ME3 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER ME2 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER ME1 ;
  RECT 0.000 109.540 1.120 112.780 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER ME4 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER ME3 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER ME2 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER ME1 ;
  RECT 0.000 101.700 1.120 104.940 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER ME4 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER ME3 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER ME2 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER ME1 ;
  RECT 0.000 93.860 1.120 97.100 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER ME4 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER ME3 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER ME2 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER ME1 ;
  RECT 0.000 86.020 1.120 89.260 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER ME4 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER ME3 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER ME2 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER ME1 ;
  RECT 0.000 46.820 1.120 50.060 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER ME4 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER ME3 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER ME2 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER ME1 ;
  RECT 0.000 38.980 1.120 42.220 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER ME4 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER ME3 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER ME2 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER ME1 ;
  RECT 0.000 31.140 1.120 34.380 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER ME4 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER ME3 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER ME2 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER ME1 ;
  RECT 0.000 23.300 1.120 26.540 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER ME4 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER ME3 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER ME2 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER ME1 ;
  RECT 0.000 15.460 1.120 18.700 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER ME4 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER ME3 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER ME2 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER ME1 ;
  RECT 0.000 7.620 1.120 10.860 ;
 END
 PORT
  LAYER ME5 ;
  RECT 517.480 348.880 521.020 350.000 ;
  LAYER ME4 ;
  RECT 517.480 348.880 521.020 350.000 ;
  LAYER ME3 ;
  RECT 517.480 348.880 521.020 350.000 ;
  LAYER ME2 ;
  RECT 517.480 348.880 521.020 350.000 ;
  LAYER ME1 ;
  RECT 517.480 348.880 521.020 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 508.800 348.880 512.340 350.000 ;
  LAYER ME4 ;
  RECT 508.800 348.880 512.340 350.000 ;
  LAYER ME3 ;
  RECT 508.800 348.880 512.340 350.000 ;
  LAYER ME2 ;
  RECT 508.800 348.880 512.340 350.000 ;
  LAYER ME1 ;
  RECT 508.800 348.880 512.340 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 500.120 348.880 503.660 350.000 ;
  LAYER ME4 ;
  RECT 500.120 348.880 503.660 350.000 ;
  LAYER ME3 ;
  RECT 500.120 348.880 503.660 350.000 ;
  LAYER ME2 ;
  RECT 500.120 348.880 503.660 350.000 ;
  LAYER ME1 ;
  RECT 500.120 348.880 503.660 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 491.440 348.880 494.980 350.000 ;
  LAYER ME4 ;
  RECT 491.440 348.880 494.980 350.000 ;
  LAYER ME3 ;
  RECT 491.440 348.880 494.980 350.000 ;
  LAYER ME2 ;
  RECT 491.440 348.880 494.980 350.000 ;
  LAYER ME1 ;
  RECT 491.440 348.880 494.980 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 482.760 348.880 486.300 350.000 ;
  LAYER ME4 ;
  RECT 482.760 348.880 486.300 350.000 ;
  LAYER ME3 ;
  RECT 482.760 348.880 486.300 350.000 ;
  LAYER ME2 ;
  RECT 482.760 348.880 486.300 350.000 ;
  LAYER ME1 ;
  RECT 482.760 348.880 486.300 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 474.080 348.880 477.620 350.000 ;
  LAYER ME4 ;
  RECT 474.080 348.880 477.620 350.000 ;
  LAYER ME3 ;
  RECT 474.080 348.880 477.620 350.000 ;
  LAYER ME2 ;
  RECT 474.080 348.880 477.620 350.000 ;
  LAYER ME1 ;
  RECT 474.080 348.880 477.620 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 413.940 348.880 417.480 350.000 ;
  LAYER ME4 ;
  RECT 413.940 348.880 417.480 350.000 ;
  LAYER ME3 ;
  RECT 413.940 348.880 417.480 350.000 ;
  LAYER ME2 ;
  RECT 413.940 348.880 417.480 350.000 ;
  LAYER ME1 ;
  RECT 413.940 348.880 417.480 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 405.260 348.880 408.800 350.000 ;
  LAYER ME4 ;
  RECT 405.260 348.880 408.800 350.000 ;
  LAYER ME3 ;
  RECT 405.260 348.880 408.800 350.000 ;
  LAYER ME2 ;
  RECT 405.260 348.880 408.800 350.000 ;
  LAYER ME1 ;
  RECT 405.260 348.880 408.800 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 396.580 348.880 400.120 350.000 ;
  LAYER ME4 ;
  RECT 396.580 348.880 400.120 350.000 ;
  LAYER ME3 ;
  RECT 396.580 348.880 400.120 350.000 ;
  LAYER ME2 ;
  RECT 396.580 348.880 400.120 350.000 ;
  LAYER ME1 ;
  RECT 396.580 348.880 400.120 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 387.900 348.880 391.440 350.000 ;
  LAYER ME4 ;
  RECT 387.900 348.880 391.440 350.000 ;
  LAYER ME3 ;
  RECT 387.900 348.880 391.440 350.000 ;
  LAYER ME2 ;
  RECT 387.900 348.880 391.440 350.000 ;
  LAYER ME1 ;
  RECT 387.900 348.880 391.440 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 379.220 348.880 382.760 350.000 ;
  LAYER ME4 ;
  RECT 379.220 348.880 382.760 350.000 ;
  LAYER ME3 ;
  RECT 379.220 348.880 382.760 350.000 ;
  LAYER ME2 ;
  RECT 379.220 348.880 382.760 350.000 ;
  LAYER ME1 ;
  RECT 379.220 348.880 382.760 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 370.540 348.880 374.080 350.000 ;
  LAYER ME4 ;
  RECT 370.540 348.880 374.080 350.000 ;
  LAYER ME3 ;
  RECT 370.540 348.880 374.080 350.000 ;
  LAYER ME2 ;
  RECT 370.540 348.880 374.080 350.000 ;
  LAYER ME1 ;
  RECT 370.540 348.880 374.080 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 310.400 348.880 313.940 350.000 ;
  LAYER ME4 ;
  RECT 310.400 348.880 313.940 350.000 ;
  LAYER ME3 ;
  RECT 310.400 348.880 313.940 350.000 ;
  LAYER ME2 ;
  RECT 310.400 348.880 313.940 350.000 ;
  LAYER ME1 ;
  RECT 310.400 348.880 313.940 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 301.720 348.880 305.260 350.000 ;
  LAYER ME4 ;
  RECT 301.720 348.880 305.260 350.000 ;
  LAYER ME3 ;
  RECT 301.720 348.880 305.260 350.000 ;
  LAYER ME2 ;
  RECT 301.720 348.880 305.260 350.000 ;
  LAYER ME1 ;
  RECT 301.720 348.880 305.260 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 255.840 348.880 259.380 350.000 ;
  LAYER ME4 ;
  RECT 255.840 348.880 259.380 350.000 ;
  LAYER ME3 ;
  RECT 255.840 348.880 259.380 350.000 ;
  LAYER ME2 ;
  RECT 255.840 348.880 259.380 350.000 ;
  LAYER ME1 ;
  RECT 255.840 348.880 259.380 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 232.900 348.880 236.440 350.000 ;
  LAYER ME4 ;
  RECT 232.900 348.880 236.440 350.000 ;
  LAYER ME3 ;
  RECT 232.900 348.880 236.440 350.000 ;
  LAYER ME2 ;
  RECT 232.900 348.880 236.440 350.000 ;
  LAYER ME1 ;
  RECT 232.900 348.880 236.440 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 224.220 348.880 227.760 350.000 ;
  LAYER ME4 ;
  RECT 224.220 348.880 227.760 350.000 ;
  LAYER ME3 ;
  RECT 224.220 348.880 227.760 350.000 ;
  LAYER ME2 ;
  RECT 224.220 348.880 227.760 350.000 ;
  LAYER ME1 ;
  RECT 224.220 348.880 227.760 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 215.540 348.880 219.080 350.000 ;
  LAYER ME4 ;
  RECT 215.540 348.880 219.080 350.000 ;
  LAYER ME3 ;
  RECT 215.540 348.880 219.080 350.000 ;
  LAYER ME2 ;
  RECT 215.540 348.880 219.080 350.000 ;
  LAYER ME1 ;
  RECT 215.540 348.880 219.080 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 172.140 348.880 175.680 350.000 ;
  LAYER ME4 ;
  RECT 172.140 348.880 175.680 350.000 ;
  LAYER ME3 ;
  RECT 172.140 348.880 175.680 350.000 ;
  LAYER ME2 ;
  RECT 172.140 348.880 175.680 350.000 ;
  LAYER ME1 ;
  RECT 172.140 348.880 175.680 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 163.460 348.880 167.000 350.000 ;
  LAYER ME4 ;
  RECT 163.460 348.880 167.000 350.000 ;
  LAYER ME3 ;
  RECT 163.460 348.880 167.000 350.000 ;
  LAYER ME2 ;
  RECT 163.460 348.880 167.000 350.000 ;
  LAYER ME1 ;
  RECT 163.460 348.880 167.000 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 149.820 348.880 153.360 350.000 ;
  LAYER ME4 ;
  RECT 149.820 348.880 153.360 350.000 ;
  LAYER ME3 ;
  RECT 149.820 348.880 153.360 350.000 ;
  LAYER ME2 ;
  RECT 149.820 348.880 153.360 350.000 ;
  LAYER ME1 ;
  RECT 149.820 348.880 153.360 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 136.180 348.880 139.720 350.000 ;
  LAYER ME4 ;
  RECT 136.180 348.880 139.720 350.000 ;
  LAYER ME3 ;
  RECT 136.180 348.880 139.720 350.000 ;
  LAYER ME2 ;
  RECT 136.180 348.880 139.720 350.000 ;
  LAYER ME1 ;
  RECT 136.180 348.880 139.720 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 123.160 348.880 126.700 350.000 ;
  LAYER ME4 ;
  RECT 123.160 348.880 126.700 350.000 ;
  LAYER ME3 ;
  RECT 123.160 348.880 126.700 350.000 ;
  LAYER ME2 ;
  RECT 123.160 348.880 126.700 350.000 ;
  LAYER ME1 ;
  RECT 123.160 348.880 126.700 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 111.380 348.880 114.920 350.000 ;
  LAYER ME4 ;
  RECT 111.380 348.880 114.920 350.000 ;
  LAYER ME3 ;
  RECT 111.380 348.880 114.920 350.000 ;
  LAYER ME2 ;
  RECT 111.380 348.880 114.920 350.000 ;
  LAYER ME1 ;
  RECT 111.380 348.880 114.920 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 67.980 348.880 71.520 350.000 ;
  LAYER ME4 ;
  RECT 67.980 348.880 71.520 350.000 ;
  LAYER ME3 ;
  RECT 67.980 348.880 71.520 350.000 ;
  LAYER ME2 ;
  RECT 67.980 348.880 71.520 350.000 ;
  LAYER ME1 ;
  RECT 67.980 348.880 71.520 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 59.300 348.880 62.840 350.000 ;
  LAYER ME4 ;
  RECT 59.300 348.880 62.840 350.000 ;
  LAYER ME3 ;
  RECT 59.300 348.880 62.840 350.000 ;
  LAYER ME2 ;
  RECT 59.300 348.880 62.840 350.000 ;
  LAYER ME1 ;
  RECT 59.300 348.880 62.840 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 46.280 348.880 49.820 350.000 ;
  LAYER ME4 ;
  RECT 46.280 348.880 49.820 350.000 ;
  LAYER ME3 ;
  RECT 46.280 348.880 49.820 350.000 ;
  LAYER ME2 ;
  RECT 46.280 348.880 49.820 350.000 ;
  LAYER ME1 ;
  RECT 46.280 348.880 49.820 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 32.640 348.880 36.180 350.000 ;
  LAYER ME4 ;
  RECT 32.640 348.880 36.180 350.000 ;
  LAYER ME3 ;
  RECT 32.640 348.880 36.180 350.000 ;
  LAYER ME2 ;
  RECT 32.640 348.880 36.180 350.000 ;
  LAYER ME1 ;
  RECT 32.640 348.880 36.180 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 19.000 348.880 22.540 350.000 ;
  LAYER ME4 ;
  RECT 19.000 348.880 22.540 350.000 ;
  LAYER ME3 ;
  RECT 19.000 348.880 22.540 350.000 ;
  LAYER ME2 ;
  RECT 19.000 348.880 22.540 350.000 ;
  LAYER ME1 ;
  RECT 19.000 348.880 22.540 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 7.220 348.880 10.760 350.000 ;
  LAYER ME4 ;
  RECT 7.220 348.880 10.760 350.000 ;
  LAYER ME3 ;
  RECT 7.220 348.880 10.760 350.000 ;
  LAYER ME2 ;
  RECT 7.220 348.880 10.760 350.000 ;
  LAYER ME1 ;
  RECT 7.220 348.880 10.760 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 517.480 0.000 521.020 1.120 ;
  LAYER ME4 ;
  RECT 517.480 0.000 521.020 1.120 ;
  LAYER ME3 ;
  RECT 517.480 0.000 521.020 1.120 ;
  LAYER ME2 ;
  RECT 517.480 0.000 521.020 1.120 ;
  LAYER ME1 ;
  RECT 517.480 0.000 521.020 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 508.800 0.000 512.340 1.120 ;
  LAYER ME4 ;
  RECT 508.800 0.000 512.340 1.120 ;
  LAYER ME3 ;
  RECT 508.800 0.000 512.340 1.120 ;
  LAYER ME2 ;
  RECT 508.800 0.000 512.340 1.120 ;
  LAYER ME1 ;
  RECT 508.800 0.000 512.340 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 500.120 0.000 503.660 1.120 ;
  LAYER ME4 ;
  RECT 500.120 0.000 503.660 1.120 ;
  LAYER ME3 ;
  RECT 500.120 0.000 503.660 1.120 ;
  LAYER ME2 ;
  RECT 500.120 0.000 503.660 1.120 ;
  LAYER ME1 ;
  RECT 500.120 0.000 503.660 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 491.440 0.000 494.980 1.120 ;
  LAYER ME4 ;
  RECT 491.440 0.000 494.980 1.120 ;
  LAYER ME3 ;
  RECT 491.440 0.000 494.980 1.120 ;
  LAYER ME2 ;
  RECT 491.440 0.000 494.980 1.120 ;
  LAYER ME1 ;
  RECT 491.440 0.000 494.980 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 482.760 0.000 486.300 1.120 ;
  LAYER ME4 ;
  RECT 482.760 0.000 486.300 1.120 ;
  LAYER ME3 ;
  RECT 482.760 0.000 486.300 1.120 ;
  LAYER ME2 ;
  RECT 482.760 0.000 486.300 1.120 ;
  LAYER ME1 ;
  RECT 482.760 0.000 486.300 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 474.080 0.000 477.620 1.120 ;
  LAYER ME4 ;
  RECT 474.080 0.000 477.620 1.120 ;
  LAYER ME3 ;
  RECT 474.080 0.000 477.620 1.120 ;
  LAYER ME2 ;
  RECT 474.080 0.000 477.620 1.120 ;
  LAYER ME1 ;
  RECT 474.080 0.000 477.620 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 413.940 0.000 417.480 1.120 ;
  LAYER ME4 ;
  RECT 413.940 0.000 417.480 1.120 ;
  LAYER ME3 ;
  RECT 413.940 0.000 417.480 1.120 ;
  LAYER ME2 ;
  RECT 413.940 0.000 417.480 1.120 ;
  LAYER ME1 ;
  RECT 413.940 0.000 417.480 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 405.260 0.000 408.800 1.120 ;
  LAYER ME4 ;
  RECT 405.260 0.000 408.800 1.120 ;
  LAYER ME3 ;
  RECT 405.260 0.000 408.800 1.120 ;
  LAYER ME2 ;
  RECT 405.260 0.000 408.800 1.120 ;
  LAYER ME1 ;
  RECT 405.260 0.000 408.800 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 396.580 0.000 400.120 1.120 ;
  LAYER ME4 ;
  RECT 396.580 0.000 400.120 1.120 ;
  LAYER ME3 ;
  RECT 396.580 0.000 400.120 1.120 ;
  LAYER ME2 ;
  RECT 396.580 0.000 400.120 1.120 ;
  LAYER ME1 ;
  RECT 396.580 0.000 400.120 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 387.900 0.000 391.440 1.120 ;
  LAYER ME4 ;
  RECT 387.900 0.000 391.440 1.120 ;
  LAYER ME3 ;
  RECT 387.900 0.000 391.440 1.120 ;
  LAYER ME2 ;
  RECT 387.900 0.000 391.440 1.120 ;
  LAYER ME1 ;
  RECT 387.900 0.000 391.440 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 379.220 0.000 382.760 1.120 ;
  LAYER ME4 ;
  RECT 379.220 0.000 382.760 1.120 ;
  LAYER ME3 ;
  RECT 379.220 0.000 382.760 1.120 ;
  LAYER ME2 ;
  RECT 379.220 0.000 382.760 1.120 ;
  LAYER ME1 ;
  RECT 379.220 0.000 382.760 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 370.540 0.000 374.080 1.120 ;
  LAYER ME4 ;
  RECT 370.540 0.000 374.080 1.120 ;
  LAYER ME3 ;
  RECT 370.540 0.000 374.080 1.120 ;
  LAYER ME2 ;
  RECT 370.540 0.000 374.080 1.120 ;
  LAYER ME1 ;
  RECT 370.540 0.000 374.080 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER ME4 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER ME3 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER ME2 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER ME1 ;
  RECT 310.400 0.000 313.940 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER ME4 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER ME3 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER ME2 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER ME1 ;
  RECT 301.720 0.000 305.260 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 255.840 0.000 259.380 1.120 ;
  LAYER ME4 ;
  RECT 255.840 0.000 259.380 1.120 ;
  LAYER ME3 ;
  RECT 255.840 0.000 259.380 1.120 ;
  LAYER ME2 ;
  RECT 255.840 0.000 259.380 1.120 ;
  LAYER ME1 ;
  RECT 255.840 0.000 259.380 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 232.900 0.000 236.440 1.120 ;
  LAYER ME4 ;
  RECT 232.900 0.000 236.440 1.120 ;
  LAYER ME3 ;
  RECT 232.900 0.000 236.440 1.120 ;
  LAYER ME2 ;
  RECT 232.900 0.000 236.440 1.120 ;
  LAYER ME1 ;
  RECT 232.900 0.000 236.440 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 224.220 0.000 227.760 1.120 ;
  LAYER ME4 ;
  RECT 224.220 0.000 227.760 1.120 ;
  LAYER ME3 ;
  RECT 224.220 0.000 227.760 1.120 ;
  LAYER ME2 ;
  RECT 224.220 0.000 227.760 1.120 ;
  LAYER ME1 ;
  RECT 224.220 0.000 227.760 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 215.540 0.000 219.080 1.120 ;
  LAYER ME4 ;
  RECT 215.540 0.000 219.080 1.120 ;
  LAYER ME3 ;
  RECT 215.540 0.000 219.080 1.120 ;
  LAYER ME2 ;
  RECT 215.540 0.000 219.080 1.120 ;
  LAYER ME1 ;
  RECT 215.540 0.000 219.080 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 172.140 0.000 175.680 1.120 ;
  LAYER ME4 ;
  RECT 172.140 0.000 175.680 1.120 ;
  LAYER ME3 ;
  RECT 172.140 0.000 175.680 1.120 ;
  LAYER ME2 ;
  RECT 172.140 0.000 175.680 1.120 ;
  LAYER ME1 ;
  RECT 172.140 0.000 175.680 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 163.460 0.000 167.000 1.120 ;
  LAYER ME4 ;
  RECT 163.460 0.000 167.000 1.120 ;
  LAYER ME3 ;
  RECT 163.460 0.000 167.000 1.120 ;
  LAYER ME2 ;
  RECT 163.460 0.000 167.000 1.120 ;
  LAYER ME1 ;
  RECT 163.460 0.000 167.000 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 149.820 0.000 153.360 1.120 ;
  LAYER ME4 ;
  RECT 149.820 0.000 153.360 1.120 ;
  LAYER ME3 ;
  RECT 149.820 0.000 153.360 1.120 ;
  LAYER ME2 ;
  RECT 149.820 0.000 153.360 1.120 ;
  LAYER ME1 ;
  RECT 149.820 0.000 153.360 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 136.180 0.000 139.720 1.120 ;
  LAYER ME4 ;
  RECT 136.180 0.000 139.720 1.120 ;
  LAYER ME3 ;
  RECT 136.180 0.000 139.720 1.120 ;
  LAYER ME2 ;
  RECT 136.180 0.000 139.720 1.120 ;
  LAYER ME1 ;
  RECT 136.180 0.000 139.720 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 123.160 0.000 126.700 1.120 ;
  LAYER ME4 ;
  RECT 123.160 0.000 126.700 1.120 ;
  LAYER ME3 ;
  RECT 123.160 0.000 126.700 1.120 ;
  LAYER ME2 ;
  RECT 123.160 0.000 126.700 1.120 ;
  LAYER ME1 ;
  RECT 123.160 0.000 126.700 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 111.380 0.000 114.920 1.120 ;
  LAYER ME4 ;
  RECT 111.380 0.000 114.920 1.120 ;
  LAYER ME3 ;
  RECT 111.380 0.000 114.920 1.120 ;
  LAYER ME2 ;
  RECT 111.380 0.000 114.920 1.120 ;
  LAYER ME1 ;
  RECT 111.380 0.000 114.920 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 67.980 0.000 71.520 1.120 ;
  LAYER ME4 ;
  RECT 67.980 0.000 71.520 1.120 ;
  LAYER ME3 ;
  RECT 67.980 0.000 71.520 1.120 ;
  LAYER ME2 ;
  RECT 67.980 0.000 71.520 1.120 ;
  LAYER ME1 ;
  RECT 67.980 0.000 71.520 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER ME4 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER ME3 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER ME2 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER ME1 ;
  RECT 59.300 0.000 62.840 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER ME4 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER ME3 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER ME2 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER ME1 ;
  RECT 46.280 0.000 49.820 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER ME4 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER ME3 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER ME2 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER ME1 ;
  RECT 32.640 0.000 36.180 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER ME4 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER ME3 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER ME2 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER ME1 ;
  RECT 19.000 0.000 22.540 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER ME4 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER ME3 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER ME2 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER ME1 ;
  RECT 7.220 0.000 10.760 1.120 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME5 ;
  RECT 543.860 332.980 544.980 336.220 ;
  LAYER ME4 ;
  RECT 543.860 332.980 544.980 336.220 ;
  LAYER ME3 ;
  RECT 543.860 332.980 544.980 336.220 ;
  LAYER ME2 ;
  RECT 543.860 332.980 544.980 336.220 ;
  LAYER ME1 ;
  RECT 543.860 332.980 544.980 336.220 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 325.140 544.980 328.380 ;
  LAYER ME4 ;
  RECT 543.860 325.140 544.980 328.380 ;
  LAYER ME3 ;
  RECT 543.860 325.140 544.980 328.380 ;
  LAYER ME2 ;
  RECT 543.860 325.140 544.980 328.380 ;
  LAYER ME1 ;
  RECT 543.860 325.140 544.980 328.380 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 285.940 544.980 289.180 ;
  LAYER ME4 ;
  RECT 543.860 285.940 544.980 289.180 ;
  LAYER ME3 ;
  RECT 543.860 285.940 544.980 289.180 ;
  LAYER ME2 ;
  RECT 543.860 285.940 544.980 289.180 ;
  LAYER ME1 ;
  RECT 543.860 285.940 544.980 289.180 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 278.100 544.980 281.340 ;
  LAYER ME4 ;
  RECT 543.860 278.100 544.980 281.340 ;
  LAYER ME3 ;
  RECT 543.860 278.100 544.980 281.340 ;
  LAYER ME2 ;
  RECT 543.860 278.100 544.980 281.340 ;
  LAYER ME1 ;
  RECT 543.860 278.100 544.980 281.340 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 270.260 544.980 273.500 ;
  LAYER ME4 ;
  RECT 543.860 270.260 544.980 273.500 ;
  LAYER ME3 ;
  RECT 543.860 270.260 544.980 273.500 ;
  LAYER ME2 ;
  RECT 543.860 270.260 544.980 273.500 ;
  LAYER ME1 ;
  RECT 543.860 270.260 544.980 273.500 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 262.420 544.980 265.660 ;
  LAYER ME4 ;
  RECT 543.860 262.420 544.980 265.660 ;
  LAYER ME3 ;
  RECT 543.860 262.420 544.980 265.660 ;
  LAYER ME2 ;
  RECT 543.860 262.420 544.980 265.660 ;
  LAYER ME1 ;
  RECT 543.860 262.420 544.980 265.660 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 254.580 544.980 257.820 ;
  LAYER ME4 ;
  RECT 543.860 254.580 544.980 257.820 ;
  LAYER ME3 ;
  RECT 543.860 254.580 544.980 257.820 ;
  LAYER ME2 ;
  RECT 543.860 254.580 544.980 257.820 ;
  LAYER ME1 ;
  RECT 543.860 254.580 544.980 257.820 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 246.740 544.980 249.980 ;
  LAYER ME4 ;
  RECT 543.860 246.740 544.980 249.980 ;
  LAYER ME3 ;
  RECT 543.860 246.740 544.980 249.980 ;
  LAYER ME2 ;
  RECT 543.860 246.740 544.980 249.980 ;
  LAYER ME1 ;
  RECT 543.860 246.740 544.980 249.980 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 207.540 544.980 210.780 ;
  LAYER ME4 ;
  RECT 543.860 207.540 544.980 210.780 ;
  LAYER ME3 ;
  RECT 543.860 207.540 544.980 210.780 ;
  LAYER ME2 ;
  RECT 543.860 207.540 544.980 210.780 ;
  LAYER ME1 ;
  RECT 543.860 207.540 544.980 210.780 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 199.700 544.980 202.940 ;
  LAYER ME4 ;
  RECT 543.860 199.700 544.980 202.940 ;
  LAYER ME3 ;
  RECT 543.860 199.700 544.980 202.940 ;
  LAYER ME2 ;
  RECT 543.860 199.700 544.980 202.940 ;
  LAYER ME1 ;
  RECT 543.860 199.700 544.980 202.940 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 191.860 544.980 195.100 ;
  LAYER ME4 ;
  RECT 543.860 191.860 544.980 195.100 ;
  LAYER ME3 ;
  RECT 543.860 191.860 544.980 195.100 ;
  LAYER ME2 ;
  RECT 543.860 191.860 544.980 195.100 ;
  LAYER ME1 ;
  RECT 543.860 191.860 544.980 195.100 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 184.020 544.980 187.260 ;
  LAYER ME4 ;
  RECT 543.860 184.020 544.980 187.260 ;
  LAYER ME3 ;
  RECT 543.860 184.020 544.980 187.260 ;
  LAYER ME2 ;
  RECT 543.860 184.020 544.980 187.260 ;
  LAYER ME1 ;
  RECT 543.860 184.020 544.980 187.260 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 176.180 544.980 179.420 ;
  LAYER ME4 ;
  RECT 543.860 176.180 544.980 179.420 ;
  LAYER ME3 ;
  RECT 543.860 176.180 544.980 179.420 ;
  LAYER ME2 ;
  RECT 543.860 176.180 544.980 179.420 ;
  LAYER ME1 ;
  RECT 543.860 176.180 544.980 179.420 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 168.340 544.980 171.580 ;
  LAYER ME4 ;
  RECT 543.860 168.340 544.980 171.580 ;
  LAYER ME3 ;
  RECT 543.860 168.340 544.980 171.580 ;
  LAYER ME2 ;
  RECT 543.860 168.340 544.980 171.580 ;
  LAYER ME1 ;
  RECT 543.860 168.340 544.980 171.580 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 129.140 544.980 132.380 ;
  LAYER ME4 ;
  RECT 543.860 129.140 544.980 132.380 ;
  LAYER ME3 ;
  RECT 543.860 129.140 544.980 132.380 ;
  LAYER ME2 ;
  RECT 543.860 129.140 544.980 132.380 ;
  LAYER ME1 ;
  RECT 543.860 129.140 544.980 132.380 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 121.300 544.980 124.540 ;
  LAYER ME4 ;
  RECT 543.860 121.300 544.980 124.540 ;
  LAYER ME3 ;
  RECT 543.860 121.300 544.980 124.540 ;
  LAYER ME2 ;
  RECT 543.860 121.300 544.980 124.540 ;
  LAYER ME1 ;
  RECT 543.860 121.300 544.980 124.540 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 113.460 544.980 116.700 ;
  LAYER ME4 ;
  RECT 543.860 113.460 544.980 116.700 ;
  LAYER ME3 ;
  RECT 543.860 113.460 544.980 116.700 ;
  LAYER ME2 ;
  RECT 543.860 113.460 544.980 116.700 ;
  LAYER ME1 ;
  RECT 543.860 113.460 544.980 116.700 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 105.620 544.980 108.860 ;
  LAYER ME4 ;
  RECT 543.860 105.620 544.980 108.860 ;
  LAYER ME3 ;
  RECT 543.860 105.620 544.980 108.860 ;
  LAYER ME2 ;
  RECT 543.860 105.620 544.980 108.860 ;
  LAYER ME1 ;
  RECT 543.860 105.620 544.980 108.860 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 97.780 544.980 101.020 ;
  LAYER ME4 ;
  RECT 543.860 97.780 544.980 101.020 ;
  LAYER ME3 ;
  RECT 543.860 97.780 544.980 101.020 ;
  LAYER ME2 ;
  RECT 543.860 97.780 544.980 101.020 ;
  LAYER ME1 ;
  RECT 543.860 97.780 544.980 101.020 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 89.940 544.980 93.180 ;
  LAYER ME4 ;
  RECT 543.860 89.940 544.980 93.180 ;
  LAYER ME3 ;
  RECT 543.860 89.940 544.980 93.180 ;
  LAYER ME2 ;
  RECT 543.860 89.940 544.980 93.180 ;
  LAYER ME1 ;
  RECT 543.860 89.940 544.980 93.180 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 50.740 544.980 53.980 ;
  LAYER ME4 ;
  RECT 543.860 50.740 544.980 53.980 ;
  LAYER ME3 ;
  RECT 543.860 50.740 544.980 53.980 ;
  LAYER ME2 ;
  RECT 543.860 50.740 544.980 53.980 ;
  LAYER ME1 ;
  RECT 543.860 50.740 544.980 53.980 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 42.900 544.980 46.140 ;
  LAYER ME4 ;
  RECT 543.860 42.900 544.980 46.140 ;
  LAYER ME3 ;
  RECT 543.860 42.900 544.980 46.140 ;
  LAYER ME2 ;
  RECT 543.860 42.900 544.980 46.140 ;
  LAYER ME1 ;
  RECT 543.860 42.900 544.980 46.140 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 35.060 544.980 38.300 ;
  LAYER ME4 ;
  RECT 543.860 35.060 544.980 38.300 ;
  LAYER ME3 ;
  RECT 543.860 35.060 544.980 38.300 ;
  LAYER ME2 ;
  RECT 543.860 35.060 544.980 38.300 ;
  LAYER ME1 ;
  RECT 543.860 35.060 544.980 38.300 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 27.220 544.980 30.460 ;
  LAYER ME4 ;
  RECT 543.860 27.220 544.980 30.460 ;
  LAYER ME3 ;
  RECT 543.860 27.220 544.980 30.460 ;
  LAYER ME2 ;
  RECT 543.860 27.220 544.980 30.460 ;
  LAYER ME1 ;
  RECT 543.860 27.220 544.980 30.460 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 19.380 544.980 22.620 ;
  LAYER ME4 ;
  RECT 543.860 19.380 544.980 22.620 ;
  LAYER ME3 ;
  RECT 543.860 19.380 544.980 22.620 ;
  LAYER ME2 ;
  RECT 543.860 19.380 544.980 22.620 ;
  LAYER ME1 ;
  RECT 543.860 19.380 544.980 22.620 ;
 END
 PORT
  LAYER ME5 ;
  RECT 543.860 11.540 544.980 14.780 ;
  LAYER ME4 ;
  RECT 543.860 11.540 544.980 14.780 ;
  LAYER ME3 ;
  RECT 543.860 11.540 544.980 14.780 ;
  LAYER ME2 ;
  RECT 543.860 11.540 544.980 14.780 ;
  LAYER ME1 ;
  RECT 543.860 11.540 544.980 14.780 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER ME4 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER ME3 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER ME2 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER ME1 ;
  RECT 0.000 332.980 1.120 336.220 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER ME4 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER ME3 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER ME2 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER ME1 ;
  RECT 0.000 325.140 1.120 328.380 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER ME4 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER ME3 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER ME2 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER ME1 ;
  RECT 0.000 285.940 1.120 289.180 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER ME4 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER ME3 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER ME2 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER ME1 ;
  RECT 0.000 278.100 1.120 281.340 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER ME4 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER ME3 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER ME2 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER ME1 ;
  RECT 0.000 270.260 1.120 273.500 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER ME4 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER ME3 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER ME2 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER ME1 ;
  RECT 0.000 262.420 1.120 265.660 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER ME4 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER ME3 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER ME2 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER ME1 ;
  RECT 0.000 254.580 1.120 257.820 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER ME4 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER ME3 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER ME2 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER ME1 ;
  RECT 0.000 246.740 1.120 249.980 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER ME4 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER ME3 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER ME2 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER ME1 ;
  RECT 0.000 207.540 1.120 210.780 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER ME4 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER ME3 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER ME2 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER ME1 ;
  RECT 0.000 199.700 1.120 202.940 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER ME4 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER ME3 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER ME2 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER ME1 ;
  RECT 0.000 191.860 1.120 195.100 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER ME4 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER ME3 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER ME2 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER ME1 ;
  RECT 0.000 184.020 1.120 187.260 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER ME4 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER ME3 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER ME2 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER ME1 ;
  RECT 0.000 176.180 1.120 179.420 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER ME4 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER ME3 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER ME2 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER ME1 ;
  RECT 0.000 168.340 1.120 171.580 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER ME4 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER ME3 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER ME2 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER ME1 ;
  RECT 0.000 129.140 1.120 132.380 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER ME4 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER ME3 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER ME2 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER ME1 ;
  RECT 0.000 121.300 1.120 124.540 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER ME4 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER ME3 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER ME2 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER ME1 ;
  RECT 0.000 113.460 1.120 116.700 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER ME4 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER ME3 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER ME2 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER ME1 ;
  RECT 0.000 105.620 1.120 108.860 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER ME4 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER ME3 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER ME2 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER ME1 ;
  RECT 0.000 97.780 1.120 101.020 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER ME4 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER ME3 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER ME2 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER ME1 ;
  RECT 0.000 89.940 1.120 93.180 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER ME4 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER ME3 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER ME2 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER ME1 ;
  RECT 0.000 50.740 1.120 53.980 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER ME4 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER ME3 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER ME2 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER ME1 ;
  RECT 0.000 42.900 1.120 46.140 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER ME4 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER ME3 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER ME2 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER ME1 ;
  RECT 0.000 35.060 1.120 38.300 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER ME4 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER ME3 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER ME2 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER ME1 ;
  RECT 0.000 27.220 1.120 30.460 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER ME4 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER ME3 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER ME2 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER ME1 ;
  RECT 0.000 19.380 1.120 22.620 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER ME4 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER ME3 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER ME2 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER ME1 ;
  RECT 0.000 11.540 1.120 14.780 ;
 END
 PORT
  LAYER ME5 ;
  RECT 521.820 348.880 525.360 350.000 ;
  LAYER ME4 ;
  RECT 521.820 348.880 525.360 350.000 ;
  LAYER ME3 ;
  RECT 521.820 348.880 525.360 350.000 ;
  LAYER ME2 ;
  RECT 521.820 348.880 525.360 350.000 ;
  LAYER ME1 ;
  RECT 521.820 348.880 525.360 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 513.140 348.880 516.680 350.000 ;
  LAYER ME4 ;
  RECT 513.140 348.880 516.680 350.000 ;
  LAYER ME3 ;
  RECT 513.140 348.880 516.680 350.000 ;
  LAYER ME2 ;
  RECT 513.140 348.880 516.680 350.000 ;
  LAYER ME1 ;
  RECT 513.140 348.880 516.680 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 504.460 348.880 508.000 350.000 ;
  LAYER ME4 ;
  RECT 504.460 348.880 508.000 350.000 ;
  LAYER ME3 ;
  RECT 504.460 348.880 508.000 350.000 ;
  LAYER ME2 ;
  RECT 504.460 348.880 508.000 350.000 ;
  LAYER ME1 ;
  RECT 504.460 348.880 508.000 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 495.780 348.880 499.320 350.000 ;
  LAYER ME4 ;
  RECT 495.780 348.880 499.320 350.000 ;
  LAYER ME3 ;
  RECT 495.780 348.880 499.320 350.000 ;
  LAYER ME2 ;
  RECT 495.780 348.880 499.320 350.000 ;
  LAYER ME1 ;
  RECT 495.780 348.880 499.320 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 487.100 348.880 490.640 350.000 ;
  LAYER ME4 ;
  RECT 487.100 348.880 490.640 350.000 ;
  LAYER ME3 ;
  RECT 487.100 348.880 490.640 350.000 ;
  LAYER ME2 ;
  RECT 487.100 348.880 490.640 350.000 ;
  LAYER ME1 ;
  RECT 487.100 348.880 490.640 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 478.420 348.880 481.960 350.000 ;
  LAYER ME4 ;
  RECT 478.420 348.880 481.960 350.000 ;
  LAYER ME3 ;
  RECT 478.420 348.880 481.960 350.000 ;
  LAYER ME2 ;
  RECT 478.420 348.880 481.960 350.000 ;
  LAYER ME1 ;
  RECT 478.420 348.880 481.960 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 418.280 348.880 421.820 350.000 ;
  LAYER ME4 ;
  RECT 418.280 348.880 421.820 350.000 ;
  LAYER ME3 ;
  RECT 418.280 348.880 421.820 350.000 ;
  LAYER ME2 ;
  RECT 418.280 348.880 421.820 350.000 ;
  LAYER ME1 ;
  RECT 418.280 348.880 421.820 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 409.600 348.880 413.140 350.000 ;
  LAYER ME4 ;
  RECT 409.600 348.880 413.140 350.000 ;
  LAYER ME3 ;
  RECT 409.600 348.880 413.140 350.000 ;
  LAYER ME2 ;
  RECT 409.600 348.880 413.140 350.000 ;
  LAYER ME1 ;
  RECT 409.600 348.880 413.140 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 400.920 348.880 404.460 350.000 ;
  LAYER ME4 ;
  RECT 400.920 348.880 404.460 350.000 ;
  LAYER ME3 ;
  RECT 400.920 348.880 404.460 350.000 ;
  LAYER ME2 ;
  RECT 400.920 348.880 404.460 350.000 ;
  LAYER ME1 ;
  RECT 400.920 348.880 404.460 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 392.240 348.880 395.780 350.000 ;
  LAYER ME4 ;
  RECT 392.240 348.880 395.780 350.000 ;
  LAYER ME3 ;
  RECT 392.240 348.880 395.780 350.000 ;
  LAYER ME2 ;
  RECT 392.240 348.880 395.780 350.000 ;
  LAYER ME1 ;
  RECT 392.240 348.880 395.780 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 383.560 348.880 387.100 350.000 ;
  LAYER ME4 ;
  RECT 383.560 348.880 387.100 350.000 ;
  LAYER ME3 ;
  RECT 383.560 348.880 387.100 350.000 ;
  LAYER ME2 ;
  RECT 383.560 348.880 387.100 350.000 ;
  LAYER ME1 ;
  RECT 383.560 348.880 387.100 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 374.880 348.880 378.420 350.000 ;
  LAYER ME4 ;
  RECT 374.880 348.880 378.420 350.000 ;
  LAYER ME3 ;
  RECT 374.880 348.880 378.420 350.000 ;
  LAYER ME2 ;
  RECT 374.880 348.880 378.420 350.000 ;
  LAYER ME1 ;
  RECT 374.880 348.880 378.420 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 314.740 348.880 318.280 350.000 ;
  LAYER ME4 ;
  RECT 314.740 348.880 318.280 350.000 ;
  LAYER ME3 ;
  RECT 314.740 348.880 318.280 350.000 ;
  LAYER ME2 ;
  RECT 314.740 348.880 318.280 350.000 ;
  LAYER ME1 ;
  RECT 314.740 348.880 318.280 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 306.060 348.880 309.600 350.000 ;
  LAYER ME4 ;
  RECT 306.060 348.880 309.600 350.000 ;
  LAYER ME3 ;
  RECT 306.060 348.880 309.600 350.000 ;
  LAYER ME2 ;
  RECT 306.060 348.880 309.600 350.000 ;
  LAYER ME1 ;
  RECT 306.060 348.880 309.600 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 275.680 348.880 279.220 350.000 ;
  LAYER ME4 ;
  RECT 275.680 348.880 279.220 350.000 ;
  LAYER ME3 ;
  RECT 275.680 348.880 279.220 350.000 ;
  LAYER ME2 ;
  RECT 275.680 348.880 279.220 350.000 ;
  LAYER ME1 ;
  RECT 275.680 348.880 279.220 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 251.500 348.880 255.040 350.000 ;
  LAYER ME4 ;
  RECT 251.500 348.880 255.040 350.000 ;
  LAYER ME3 ;
  RECT 251.500 348.880 255.040 350.000 ;
  LAYER ME2 ;
  RECT 251.500 348.880 255.040 350.000 ;
  LAYER ME1 ;
  RECT 251.500 348.880 255.040 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 228.560 348.880 232.100 350.000 ;
  LAYER ME4 ;
  RECT 228.560 348.880 232.100 350.000 ;
  LAYER ME3 ;
  RECT 228.560 348.880 232.100 350.000 ;
  LAYER ME2 ;
  RECT 228.560 348.880 232.100 350.000 ;
  LAYER ME1 ;
  RECT 228.560 348.880 232.100 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 219.880 348.880 223.420 350.000 ;
  LAYER ME4 ;
  RECT 219.880 348.880 223.420 350.000 ;
  LAYER ME3 ;
  RECT 219.880 348.880 223.420 350.000 ;
  LAYER ME2 ;
  RECT 219.880 348.880 223.420 350.000 ;
  LAYER ME1 ;
  RECT 219.880 348.880 223.420 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 176.480 348.880 180.020 350.000 ;
  LAYER ME4 ;
  RECT 176.480 348.880 180.020 350.000 ;
  LAYER ME3 ;
  RECT 176.480 348.880 180.020 350.000 ;
  LAYER ME2 ;
  RECT 176.480 348.880 180.020 350.000 ;
  LAYER ME1 ;
  RECT 176.480 348.880 180.020 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 167.800 348.880 171.340 350.000 ;
  LAYER ME4 ;
  RECT 167.800 348.880 171.340 350.000 ;
  LAYER ME3 ;
  RECT 167.800 348.880 171.340 350.000 ;
  LAYER ME2 ;
  RECT 167.800 348.880 171.340 350.000 ;
  LAYER ME1 ;
  RECT 167.800 348.880 171.340 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 154.160 348.880 157.700 350.000 ;
  LAYER ME4 ;
  RECT 154.160 348.880 157.700 350.000 ;
  LAYER ME3 ;
  RECT 154.160 348.880 157.700 350.000 ;
  LAYER ME2 ;
  RECT 154.160 348.880 157.700 350.000 ;
  LAYER ME1 ;
  RECT 154.160 348.880 157.700 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 140.520 348.880 144.060 350.000 ;
  LAYER ME4 ;
  RECT 140.520 348.880 144.060 350.000 ;
  LAYER ME3 ;
  RECT 140.520 348.880 144.060 350.000 ;
  LAYER ME2 ;
  RECT 140.520 348.880 144.060 350.000 ;
  LAYER ME1 ;
  RECT 140.520 348.880 144.060 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 127.500 348.880 131.040 350.000 ;
  LAYER ME4 ;
  RECT 127.500 348.880 131.040 350.000 ;
  LAYER ME3 ;
  RECT 127.500 348.880 131.040 350.000 ;
  LAYER ME2 ;
  RECT 127.500 348.880 131.040 350.000 ;
  LAYER ME1 ;
  RECT 127.500 348.880 131.040 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 115.720 348.880 119.260 350.000 ;
  LAYER ME4 ;
  RECT 115.720 348.880 119.260 350.000 ;
  LAYER ME3 ;
  RECT 115.720 348.880 119.260 350.000 ;
  LAYER ME2 ;
  RECT 115.720 348.880 119.260 350.000 ;
  LAYER ME1 ;
  RECT 115.720 348.880 119.260 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 72.320 348.880 75.860 350.000 ;
  LAYER ME4 ;
  RECT 72.320 348.880 75.860 350.000 ;
  LAYER ME3 ;
  RECT 72.320 348.880 75.860 350.000 ;
  LAYER ME2 ;
  RECT 72.320 348.880 75.860 350.000 ;
  LAYER ME1 ;
  RECT 72.320 348.880 75.860 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 63.640 348.880 67.180 350.000 ;
  LAYER ME4 ;
  RECT 63.640 348.880 67.180 350.000 ;
  LAYER ME3 ;
  RECT 63.640 348.880 67.180 350.000 ;
  LAYER ME2 ;
  RECT 63.640 348.880 67.180 350.000 ;
  LAYER ME1 ;
  RECT 63.640 348.880 67.180 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 54.960 348.880 58.500 350.000 ;
  LAYER ME4 ;
  RECT 54.960 348.880 58.500 350.000 ;
  LAYER ME3 ;
  RECT 54.960 348.880 58.500 350.000 ;
  LAYER ME2 ;
  RECT 54.960 348.880 58.500 350.000 ;
  LAYER ME1 ;
  RECT 54.960 348.880 58.500 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 41.940 348.880 45.480 350.000 ;
  LAYER ME4 ;
  RECT 41.940 348.880 45.480 350.000 ;
  LAYER ME3 ;
  RECT 41.940 348.880 45.480 350.000 ;
  LAYER ME2 ;
  RECT 41.940 348.880 45.480 350.000 ;
  LAYER ME1 ;
  RECT 41.940 348.880 45.480 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 28.300 348.880 31.840 350.000 ;
  LAYER ME4 ;
  RECT 28.300 348.880 31.840 350.000 ;
  LAYER ME3 ;
  RECT 28.300 348.880 31.840 350.000 ;
  LAYER ME2 ;
  RECT 28.300 348.880 31.840 350.000 ;
  LAYER ME1 ;
  RECT 28.300 348.880 31.840 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 14.660 348.880 18.200 350.000 ;
  LAYER ME4 ;
  RECT 14.660 348.880 18.200 350.000 ;
  LAYER ME3 ;
  RECT 14.660 348.880 18.200 350.000 ;
  LAYER ME2 ;
  RECT 14.660 348.880 18.200 350.000 ;
  LAYER ME1 ;
  RECT 14.660 348.880 18.200 350.000 ;
 END
 PORT
  LAYER ME5 ;
  RECT 521.820 0.000 525.360 1.120 ;
  LAYER ME4 ;
  RECT 521.820 0.000 525.360 1.120 ;
  LAYER ME3 ;
  RECT 521.820 0.000 525.360 1.120 ;
  LAYER ME2 ;
  RECT 521.820 0.000 525.360 1.120 ;
  LAYER ME1 ;
  RECT 521.820 0.000 525.360 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 513.140 0.000 516.680 1.120 ;
  LAYER ME4 ;
  RECT 513.140 0.000 516.680 1.120 ;
  LAYER ME3 ;
  RECT 513.140 0.000 516.680 1.120 ;
  LAYER ME2 ;
  RECT 513.140 0.000 516.680 1.120 ;
  LAYER ME1 ;
  RECT 513.140 0.000 516.680 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 504.460 0.000 508.000 1.120 ;
  LAYER ME4 ;
  RECT 504.460 0.000 508.000 1.120 ;
  LAYER ME3 ;
  RECT 504.460 0.000 508.000 1.120 ;
  LAYER ME2 ;
  RECT 504.460 0.000 508.000 1.120 ;
  LAYER ME1 ;
  RECT 504.460 0.000 508.000 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 495.780 0.000 499.320 1.120 ;
  LAYER ME4 ;
  RECT 495.780 0.000 499.320 1.120 ;
  LAYER ME3 ;
  RECT 495.780 0.000 499.320 1.120 ;
  LAYER ME2 ;
  RECT 495.780 0.000 499.320 1.120 ;
  LAYER ME1 ;
  RECT 495.780 0.000 499.320 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 487.100 0.000 490.640 1.120 ;
  LAYER ME4 ;
  RECT 487.100 0.000 490.640 1.120 ;
  LAYER ME3 ;
  RECT 487.100 0.000 490.640 1.120 ;
  LAYER ME2 ;
  RECT 487.100 0.000 490.640 1.120 ;
  LAYER ME1 ;
  RECT 487.100 0.000 490.640 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 478.420 0.000 481.960 1.120 ;
  LAYER ME4 ;
  RECT 478.420 0.000 481.960 1.120 ;
  LAYER ME3 ;
  RECT 478.420 0.000 481.960 1.120 ;
  LAYER ME2 ;
  RECT 478.420 0.000 481.960 1.120 ;
  LAYER ME1 ;
  RECT 478.420 0.000 481.960 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER ME4 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER ME3 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER ME2 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER ME1 ;
  RECT 418.280 0.000 421.820 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 409.600 0.000 413.140 1.120 ;
  LAYER ME4 ;
  RECT 409.600 0.000 413.140 1.120 ;
  LAYER ME3 ;
  RECT 409.600 0.000 413.140 1.120 ;
  LAYER ME2 ;
  RECT 409.600 0.000 413.140 1.120 ;
  LAYER ME1 ;
  RECT 409.600 0.000 413.140 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 400.920 0.000 404.460 1.120 ;
  LAYER ME4 ;
  RECT 400.920 0.000 404.460 1.120 ;
  LAYER ME3 ;
  RECT 400.920 0.000 404.460 1.120 ;
  LAYER ME2 ;
  RECT 400.920 0.000 404.460 1.120 ;
  LAYER ME1 ;
  RECT 400.920 0.000 404.460 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 392.240 0.000 395.780 1.120 ;
  LAYER ME4 ;
  RECT 392.240 0.000 395.780 1.120 ;
  LAYER ME3 ;
  RECT 392.240 0.000 395.780 1.120 ;
  LAYER ME2 ;
  RECT 392.240 0.000 395.780 1.120 ;
  LAYER ME1 ;
  RECT 392.240 0.000 395.780 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 383.560 0.000 387.100 1.120 ;
  LAYER ME4 ;
  RECT 383.560 0.000 387.100 1.120 ;
  LAYER ME3 ;
  RECT 383.560 0.000 387.100 1.120 ;
  LAYER ME2 ;
  RECT 383.560 0.000 387.100 1.120 ;
  LAYER ME1 ;
  RECT 383.560 0.000 387.100 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 374.880 0.000 378.420 1.120 ;
  LAYER ME4 ;
  RECT 374.880 0.000 378.420 1.120 ;
  LAYER ME3 ;
  RECT 374.880 0.000 378.420 1.120 ;
  LAYER ME2 ;
  RECT 374.880 0.000 378.420 1.120 ;
  LAYER ME1 ;
  RECT 374.880 0.000 378.420 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER ME4 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER ME3 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER ME2 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER ME1 ;
  RECT 314.740 0.000 318.280 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 306.060 0.000 309.600 1.120 ;
  LAYER ME4 ;
  RECT 306.060 0.000 309.600 1.120 ;
  LAYER ME3 ;
  RECT 306.060 0.000 309.600 1.120 ;
  LAYER ME2 ;
  RECT 306.060 0.000 309.600 1.120 ;
  LAYER ME1 ;
  RECT 306.060 0.000 309.600 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 275.680 0.000 279.220 1.120 ;
  LAYER ME4 ;
  RECT 275.680 0.000 279.220 1.120 ;
  LAYER ME3 ;
  RECT 275.680 0.000 279.220 1.120 ;
  LAYER ME2 ;
  RECT 275.680 0.000 279.220 1.120 ;
  LAYER ME1 ;
  RECT 275.680 0.000 279.220 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 251.500 0.000 255.040 1.120 ;
  LAYER ME4 ;
  RECT 251.500 0.000 255.040 1.120 ;
  LAYER ME3 ;
  RECT 251.500 0.000 255.040 1.120 ;
  LAYER ME2 ;
  RECT 251.500 0.000 255.040 1.120 ;
  LAYER ME1 ;
  RECT 251.500 0.000 255.040 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 228.560 0.000 232.100 1.120 ;
  LAYER ME4 ;
  RECT 228.560 0.000 232.100 1.120 ;
  LAYER ME3 ;
  RECT 228.560 0.000 232.100 1.120 ;
  LAYER ME2 ;
  RECT 228.560 0.000 232.100 1.120 ;
  LAYER ME1 ;
  RECT 228.560 0.000 232.100 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 219.880 0.000 223.420 1.120 ;
  LAYER ME4 ;
  RECT 219.880 0.000 223.420 1.120 ;
  LAYER ME3 ;
  RECT 219.880 0.000 223.420 1.120 ;
  LAYER ME2 ;
  RECT 219.880 0.000 223.420 1.120 ;
  LAYER ME1 ;
  RECT 219.880 0.000 223.420 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER ME4 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER ME3 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER ME2 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER ME1 ;
  RECT 176.480 0.000 180.020 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 167.800 0.000 171.340 1.120 ;
  LAYER ME4 ;
  RECT 167.800 0.000 171.340 1.120 ;
  LAYER ME3 ;
  RECT 167.800 0.000 171.340 1.120 ;
  LAYER ME2 ;
  RECT 167.800 0.000 171.340 1.120 ;
  LAYER ME1 ;
  RECT 167.800 0.000 171.340 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 154.160 0.000 157.700 1.120 ;
  LAYER ME4 ;
  RECT 154.160 0.000 157.700 1.120 ;
  LAYER ME3 ;
  RECT 154.160 0.000 157.700 1.120 ;
  LAYER ME2 ;
  RECT 154.160 0.000 157.700 1.120 ;
  LAYER ME1 ;
  RECT 154.160 0.000 157.700 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER ME4 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER ME3 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER ME2 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER ME1 ;
  RECT 140.520 0.000 144.060 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 127.500 0.000 131.040 1.120 ;
  LAYER ME4 ;
  RECT 127.500 0.000 131.040 1.120 ;
  LAYER ME3 ;
  RECT 127.500 0.000 131.040 1.120 ;
  LAYER ME2 ;
  RECT 127.500 0.000 131.040 1.120 ;
  LAYER ME1 ;
  RECT 127.500 0.000 131.040 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 115.720 0.000 119.260 1.120 ;
  LAYER ME4 ;
  RECT 115.720 0.000 119.260 1.120 ;
  LAYER ME3 ;
  RECT 115.720 0.000 119.260 1.120 ;
  LAYER ME2 ;
  RECT 115.720 0.000 119.260 1.120 ;
  LAYER ME1 ;
  RECT 115.720 0.000 119.260 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 72.320 0.000 75.860 1.120 ;
  LAYER ME4 ;
  RECT 72.320 0.000 75.860 1.120 ;
  LAYER ME3 ;
  RECT 72.320 0.000 75.860 1.120 ;
  LAYER ME2 ;
  RECT 72.320 0.000 75.860 1.120 ;
  LAYER ME1 ;
  RECT 72.320 0.000 75.860 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 63.640 0.000 67.180 1.120 ;
  LAYER ME4 ;
  RECT 63.640 0.000 67.180 1.120 ;
  LAYER ME3 ;
  RECT 63.640 0.000 67.180 1.120 ;
  LAYER ME2 ;
  RECT 63.640 0.000 67.180 1.120 ;
  LAYER ME1 ;
  RECT 63.640 0.000 67.180 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER ME4 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER ME3 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER ME2 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER ME1 ;
  RECT 54.960 0.000 58.500 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER ME4 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER ME3 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER ME2 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER ME1 ;
  RECT 41.940 0.000 45.480 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER ME4 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER ME3 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER ME2 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER ME1 ;
  RECT 28.300 0.000 31.840 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER ME4 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER ME3 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER ME2 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER ME1 ;
  RECT 14.660 0.000 18.200 1.120 ;
 END
END GND
PIN DIB7
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 467.540 348.880 468.660 350.000 ;
  LAYER ME4 ;
  RECT 467.540 348.880 468.660 350.000 ;
  LAYER ME3 ;
  RECT 467.540 348.880 468.660 350.000 ;
  LAYER ME2 ;
  RECT 467.540 348.880 468.660 350.000 ;
  LAYER ME1 ;
  RECT 467.540 348.880 468.660 350.000 ;
 END
END DIB7
PIN DOB7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 454.520 348.880 455.640 350.000 ;
  LAYER ME4 ;
  RECT 454.520 348.880 455.640 350.000 ;
  LAYER ME3 ;
  RECT 454.520 348.880 455.640 350.000 ;
  LAYER ME2 ;
  RECT 454.520 348.880 455.640 350.000 ;
  LAYER ME1 ;
  RECT 454.520 348.880 455.640 350.000 ;
 END
END DOB7
PIN DIB6
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 440.880 348.880 442.000 350.000 ;
  LAYER ME4 ;
  RECT 440.880 348.880 442.000 350.000 ;
  LAYER ME3 ;
  RECT 440.880 348.880 442.000 350.000 ;
  LAYER ME2 ;
  RECT 440.880 348.880 442.000 350.000 ;
  LAYER ME1 ;
  RECT 440.880 348.880 442.000 350.000 ;
 END
END DIB6
PIN DOB6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 427.240 348.880 428.360 350.000 ;
  LAYER ME4 ;
  RECT 427.240 348.880 428.360 350.000 ;
  LAYER ME3 ;
  RECT 427.240 348.880 428.360 350.000 ;
  LAYER ME2 ;
  RECT 427.240 348.880 428.360 350.000 ;
  LAYER ME1 ;
  RECT 427.240 348.880 428.360 350.000 ;
 END
END DOB6
PIN DIB5
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 359.660 348.880 360.780 350.000 ;
  LAYER ME4 ;
  RECT 359.660 348.880 360.780 350.000 ;
  LAYER ME3 ;
  RECT 359.660 348.880 360.780 350.000 ;
  LAYER ME2 ;
  RECT 359.660 348.880 360.780 350.000 ;
  LAYER ME1 ;
  RECT 359.660 348.880 360.780 350.000 ;
 END
END DIB5
PIN DOB5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 346.020 348.880 347.140 350.000 ;
  LAYER ME4 ;
  RECT 346.020 348.880 347.140 350.000 ;
  LAYER ME3 ;
  RECT 346.020 348.880 347.140 350.000 ;
  LAYER ME2 ;
  RECT 346.020 348.880 347.140 350.000 ;
  LAYER ME1 ;
  RECT 346.020 348.880 347.140 350.000 ;
 END
END DOB5
PIN DIB4
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 333.000 348.880 334.120 350.000 ;
  LAYER ME4 ;
  RECT 333.000 348.880 334.120 350.000 ;
  LAYER ME3 ;
  RECT 333.000 348.880 334.120 350.000 ;
  LAYER ME2 ;
  RECT 333.000 348.880 334.120 350.000 ;
  LAYER ME1 ;
  RECT 333.000 348.880 334.120 350.000 ;
 END
END DIB4
PIN DOB4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 319.360 348.880 320.480 350.000 ;
  LAYER ME4 ;
  RECT 319.360 348.880 320.480 350.000 ;
  LAYER ME3 ;
  RECT 319.360 348.880 320.480 350.000 ;
  LAYER ME2 ;
  RECT 319.360 348.880 320.480 350.000 ;
  LAYER ME1 ;
  RECT 319.360 348.880 320.480 350.000 ;
 END
END DOB4
PIN B3
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 299.520 348.880 300.640 350.000 ;
  LAYER ME4 ;
  RECT 299.520 348.880 300.640 350.000 ;
  LAYER ME3 ;
  RECT 299.520 348.880 300.640 350.000 ;
  LAYER ME2 ;
  RECT 299.520 348.880 300.640 350.000 ;
  LAYER ME1 ;
  RECT 299.520 348.880 300.640 350.000 ;
 END
END B3
PIN CKB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 297.660 348.880 298.780 350.000 ;
  LAYER ME4 ;
  RECT 297.660 348.880 298.780 350.000 ;
  LAYER ME3 ;
  RECT 297.660 348.880 298.780 350.000 ;
  LAYER ME2 ;
  RECT 297.660 348.880 298.780 350.000 ;
  LAYER ME1 ;
  RECT 297.660 348.880 298.780 350.000 ;
 END
END CKB
PIN CSB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 295.180 348.880 296.300 350.000 ;
  LAYER ME4 ;
  RECT 295.180 348.880 296.300 350.000 ;
  LAYER ME3 ;
  RECT 295.180 348.880 296.300 350.000 ;
  LAYER ME2 ;
  RECT 295.180 348.880 296.300 350.000 ;
  LAYER ME1 ;
  RECT 295.180 348.880 296.300 350.000 ;
 END
END CSB
PIN WEBN
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 293.320 348.880 294.440 350.000 ;
  LAYER ME4 ;
  RECT 293.320 348.880 294.440 350.000 ;
  LAYER ME3 ;
  RECT 293.320 348.880 294.440 350.000 ;
  LAYER ME2 ;
  RECT 293.320 348.880 294.440 350.000 ;
  LAYER ME1 ;
  RECT 293.320 348.880 294.440 350.000 ;
 END
END WEBN
PIN B2
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 289.600 348.880 290.720 350.000 ;
  LAYER ME4 ;
  RECT 289.600 348.880 290.720 350.000 ;
  LAYER ME3 ;
  RECT 289.600 348.880 290.720 350.000 ;
  LAYER ME2 ;
  RECT 289.600 348.880 290.720 350.000 ;
  LAYER ME1 ;
  RECT 289.600 348.880 290.720 350.000 ;
 END
END B2
PIN OEB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 285.880 348.880 287.000 350.000 ;
  LAYER ME4 ;
  RECT 285.880 348.880 287.000 350.000 ;
  LAYER ME3 ;
  RECT 285.880 348.880 287.000 350.000 ;
  LAYER ME2 ;
  RECT 285.880 348.880 287.000 350.000 ;
  LAYER ME1 ;
  RECT 285.880 348.880 287.000 350.000 ;
 END
END OEB
PIN B1
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 284.020 348.880 285.140 350.000 ;
  LAYER ME4 ;
  RECT 284.020 348.880 285.140 350.000 ;
  LAYER ME3 ;
  RECT 284.020 348.880 285.140 350.000 ;
  LAYER ME2 ;
  RECT 284.020 348.880 285.140 350.000 ;
  LAYER ME1 ;
  RECT 284.020 348.880 285.140 350.000 ;
 END
END B1
PIN B0
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 282.160 348.880 283.280 350.000 ;
  LAYER ME4 ;
  RECT 282.160 348.880 283.280 350.000 ;
  LAYER ME3 ;
  RECT 282.160 348.880 283.280 350.000 ;
  LAYER ME2 ;
  RECT 282.160 348.880 283.280 350.000 ;
  LAYER ME1 ;
  RECT 282.160 348.880 283.280 350.000 ;
 END
END B0
PIN B6
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 273.480 348.880 274.600 350.000 ;
  LAYER ME4 ;
  RECT 273.480 348.880 274.600 350.000 ;
  LAYER ME3 ;
  RECT 273.480 348.880 274.600 350.000 ;
  LAYER ME2 ;
  RECT 273.480 348.880 274.600 350.000 ;
  LAYER ME1 ;
  RECT 273.480 348.880 274.600 350.000 ;
 END
END B6
PIN B5
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 267.900 348.880 269.020 350.000 ;
  LAYER ME4 ;
  RECT 267.900 348.880 269.020 350.000 ;
  LAYER ME3 ;
  RECT 267.900 348.880 269.020 350.000 ;
  LAYER ME2 ;
  RECT 267.900 348.880 269.020 350.000 ;
  LAYER ME1 ;
  RECT 267.900 348.880 269.020 350.000 ;
 END
END B5
PIN B4
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 262.320 348.880 263.440 350.000 ;
  LAYER ME4 ;
  RECT 262.320 348.880 263.440 350.000 ;
  LAYER ME3 ;
  RECT 262.320 348.880 263.440 350.000 ;
  LAYER ME2 ;
  RECT 262.320 348.880 263.440 350.000 ;
  LAYER ME1 ;
  RECT 262.320 348.880 263.440 350.000 ;
 END
END B4
PIN B9
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 249.300 348.880 250.420 350.000 ;
  LAYER ME4 ;
  RECT 249.300 348.880 250.420 350.000 ;
  LAYER ME3 ;
  RECT 249.300 348.880 250.420 350.000 ;
  LAYER ME2 ;
  RECT 249.300 348.880 250.420 350.000 ;
  LAYER ME1 ;
  RECT 249.300 348.880 250.420 350.000 ;
 END
END B9
PIN B8
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 243.720 348.880 244.840 350.000 ;
  LAYER ME4 ;
  RECT 243.720 348.880 244.840 350.000 ;
  LAYER ME3 ;
  RECT 243.720 348.880 244.840 350.000 ;
  LAYER ME2 ;
  RECT 243.720 348.880 244.840 350.000 ;
  LAYER ME1 ;
  RECT 243.720 348.880 244.840 350.000 ;
 END
END B8
PIN B7
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 237.520 348.880 238.640 350.000 ;
  LAYER ME4 ;
  RECT 237.520 348.880 238.640 350.000 ;
  LAYER ME3 ;
  RECT 237.520 348.880 238.640 350.000 ;
  LAYER ME2 ;
  RECT 237.520 348.880 238.640 350.000 ;
  LAYER ME1 ;
  RECT 237.520 348.880 238.640 350.000 ;
 END
END B7
PIN DIB3
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 161.260 348.880 162.380 350.000 ;
  LAYER ME4 ;
  RECT 161.260 348.880 162.380 350.000 ;
  LAYER ME3 ;
  RECT 161.260 348.880 162.380 350.000 ;
  LAYER ME2 ;
  RECT 161.260 348.880 162.380 350.000 ;
  LAYER ME1 ;
  RECT 161.260 348.880 162.380 350.000 ;
 END
END DIB3
PIN DOB3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 147.620 348.880 148.740 350.000 ;
  LAYER ME4 ;
  RECT 147.620 348.880 148.740 350.000 ;
  LAYER ME3 ;
  RECT 147.620 348.880 148.740 350.000 ;
  LAYER ME2 ;
  RECT 147.620 348.880 148.740 350.000 ;
  LAYER ME1 ;
  RECT 147.620 348.880 148.740 350.000 ;
 END
END DOB3
PIN DIB2
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 133.980 348.880 135.100 350.000 ;
  LAYER ME4 ;
  RECT 133.980 348.880 135.100 350.000 ;
  LAYER ME3 ;
  RECT 133.980 348.880 135.100 350.000 ;
  LAYER ME2 ;
  RECT 133.980 348.880 135.100 350.000 ;
  LAYER ME1 ;
  RECT 133.980 348.880 135.100 350.000 ;
 END
END DIB2
PIN DOB2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 120.960 348.880 122.080 350.000 ;
  LAYER ME4 ;
  RECT 120.960 348.880 122.080 350.000 ;
  LAYER ME3 ;
  RECT 120.960 348.880 122.080 350.000 ;
  LAYER ME2 ;
  RECT 120.960 348.880 122.080 350.000 ;
  LAYER ME1 ;
  RECT 120.960 348.880 122.080 350.000 ;
 END
END DOB2
PIN DIB1
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 52.760 348.880 53.880 350.000 ;
  LAYER ME4 ;
  RECT 52.760 348.880 53.880 350.000 ;
  LAYER ME3 ;
  RECT 52.760 348.880 53.880 350.000 ;
  LAYER ME2 ;
  RECT 52.760 348.880 53.880 350.000 ;
  LAYER ME1 ;
  RECT 52.760 348.880 53.880 350.000 ;
 END
END DIB1
PIN DOB1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 39.740 348.880 40.860 350.000 ;
  LAYER ME4 ;
  RECT 39.740 348.880 40.860 350.000 ;
  LAYER ME3 ;
  RECT 39.740 348.880 40.860 350.000 ;
  LAYER ME2 ;
  RECT 39.740 348.880 40.860 350.000 ;
  LAYER ME1 ;
  RECT 39.740 348.880 40.860 350.000 ;
 END
END DOB1
PIN DIB0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 26.100 348.880 27.220 350.000 ;
  LAYER ME4 ;
  RECT 26.100 348.880 27.220 350.000 ;
  LAYER ME3 ;
  RECT 26.100 348.880 27.220 350.000 ;
  LAYER ME2 ;
  RECT 26.100 348.880 27.220 350.000 ;
  LAYER ME1 ;
  RECT 26.100 348.880 27.220 350.000 ;
 END
END DIB0
PIN DOB0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 12.460 348.880 13.580 350.000 ;
  LAYER ME4 ;
  RECT 12.460 348.880 13.580 350.000 ;
  LAYER ME3 ;
  RECT 12.460 348.880 13.580 350.000 ;
  LAYER ME2 ;
  RECT 12.460 348.880 13.580 350.000 ;
  LAYER ME1 ;
  RECT 12.460 348.880 13.580 350.000 ;
 END
END DOB0
PIN DIA7
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 467.540 0.000 468.660 1.120 ;
  LAYER ME4 ;
  RECT 467.540 0.000 468.660 1.120 ;
  LAYER ME3 ;
  RECT 467.540 0.000 468.660 1.120 ;
  LAYER ME2 ;
  RECT 467.540 0.000 468.660 1.120 ;
  LAYER ME1 ;
  RECT 467.540 0.000 468.660 1.120 ;
 END
END DIA7
PIN DOA7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 454.520 0.000 455.640 1.120 ;
  LAYER ME4 ;
  RECT 454.520 0.000 455.640 1.120 ;
  LAYER ME3 ;
  RECT 454.520 0.000 455.640 1.120 ;
  LAYER ME2 ;
  RECT 454.520 0.000 455.640 1.120 ;
  LAYER ME1 ;
  RECT 454.520 0.000 455.640 1.120 ;
 END
END DOA7
PIN DIA6
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 440.880 0.000 442.000 1.120 ;
  LAYER ME4 ;
  RECT 440.880 0.000 442.000 1.120 ;
  LAYER ME3 ;
  RECT 440.880 0.000 442.000 1.120 ;
  LAYER ME2 ;
  RECT 440.880 0.000 442.000 1.120 ;
  LAYER ME1 ;
  RECT 440.880 0.000 442.000 1.120 ;
 END
END DIA6
PIN DOA6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 427.240 0.000 428.360 1.120 ;
  LAYER ME4 ;
  RECT 427.240 0.000 428.360 1.120 ;
  LAYER ME3 ;
  RECT 427.240 0.000 428.360 1.120 ;
  LAYER ME2 ;
  RECT 427.240 0.000 428.360 1.120 ;
  LAYER ME1 ;
  RECT 427.240 0.000 428.360 1.120 ;
 END
END DOA6
PIN DIA5
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 359.660 0.000 360.780 1.120 ;
  LAYER ME4 ;
  RECT 359.660 0.000 360.780 1.120 ;
  LAYER ME3 ;
  RECT 359.660 0.000 360.780 1.120 ;
  LAYER ME2 ;
  RECT 359.660 0.000 360.780 1.120 ;
  LAYER ME1 ;
  RECT 359.660 0.000 360.780 1.120 ;
 END
END DIA5
PIN DOA5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER ME4 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER ME3 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER ME2 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER ME1 ;
  RECT 346.020 0.000 347.140 1.120 ;
 END
END DOA5
PIN DIA4
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 333.000 0.000 334.120 1.120 ;
  LAYER ME4 ;
  RECT 333.000 0.000 334.120 1.120 ;
  LAYER ME3 ;
  RECT 333.000 0.000 334.120 1.120 ;
  LAYER ME2 ;
  RECT 333.000 0.000 334.120 1.120 ;
  LAYER ME1 ;
  RECT 333.000 0.000 334.120 1.120 ;
 END
END DIA4
PIN DOA4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 319.360 0.000 320.480 1.120 ;
  LAYER ME4 ;
  RECT 319.360 0.000 320.480 1.120 ;
  LAYER ME3 ;
  RECT 319.360 0.000 320.480 1.120 ;
  LAYER ME2 ;
  RECT 319.360 0.000 320.480 1.120 ;
  LAYER ME1 ;
  RECT 319.360 0.000 320.480 1.120 ;
 END
END DOA4
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 299.520 0.000 300.640 1.120 ;
  LAYER ME4 ;
  RECT 299.520 0.000 300.640 1.120 ;
  LAYER ME3 ;
  RECT 299.520 0.000 300.640 1.120 ;
  LAYER ME2 ;
  RECT 299.520 0.000 300.640 1.120 ;
  LAYER ME1 ;
  RECT 299.520 0.000 300.640 1.120 ;
 END
END A3
PIN CKA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 297.660 0.000 298.780 1.120 ;
  LAYER ME4 ;
  RECT 297.660 0.000 298.780 1.120 ;
  LAYER ME3 ;
  RECT 297.660 0.000 298.780 1.120 ;
  LAYER ME2 ;
  RECT 297.660 0.000 298.780 1.120 ;
  LAYER ME1 ;
  RECT 297.660 0.000 298.780 1.120 ;
 END
END CKA
PIN CSA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER ME4 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER ME3 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER ME2 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER ME1 ;
  RECT 295.180 0.000 296.300 1.120 ;
 END
END CSA
PIN WEAN
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 293.320 0.000 294.440 1.120 ;
  LAYER ME4 ;
  RECT 293.320 0.000 294.440 1.120 ;
  LAYER ME3 ;
  RECT 293.320 0.000 294.440 1.120 ;
  LAYER ME2 ;
  RECT 293.320 0.000 294.440 1.120 ;
  LAYER ME1 ;
  RECT 293.320 0.000 294.440 1.120 ;
 END
END WEAN
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME4 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME3 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME2 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME1 ;
  RECT 289.600 0.000 290.720 1.120 ;
 END
END A2
PIN OEA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 285.880 0.000 287.000 1.120 ;
  LAYER ME4 ;
  RECT 285.880 0.000 287.000 1.120 ;
  LAYER ME3 ;
  RECT 285.880 0.000 287.000 1.120 ;
  LAYER ME2 ;
  RECT 285.880 0.000 287.000 1.120 ;
  LAYER ME1 ;
  RECT 285.880 0.000 287.000 1.120 ;
 END
END OEA
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 284.020 0.000 285.140 1.120 ;
  LAYER ME4 ;
  RECT 284.020 0.000 285.140 1.120 ;
  LAYER ME3 ;
  RECT 284.020 0.000 285.140 1.120 ;
  LAYER ME2 ;
  RECT 284.020 0.000 285.140 1.120 ;
  LAYER ME1 ;
  RECT 284.020 0.000 285.140 1.120 ;
 END
END A1
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 282.160 0.000 283.280 1.120 ;
  LAYER ME4 ;
  RECT 282.160 0.000 283.280 1.120 ;
  LAYER ME3 ;
  RECT 282.160 0.000 283.280 1.120 ;
  LAYER ME2 ;
  RECT 282.160 0.000 283.280 1.120 ;
  LAYER ME1 ;
  RECT 282.160 0.000 283.280 1.120 ;
 END
END A0
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 273.480 0.000 274.600 1.120 ;
  LAYER ME4 ;
  RECT 273.480 0.000 274.600 1.120 ;
  LAYER ME3 ;
  RECT 273.480 0.000 274.600 1.120 ;
  LAYER ME2 ;
  RECT 273.480 0.000 274.600 1.120 ;
  LAYER ME1 ;
  RECT 273.480 0.000 274.600 1.120 ;
 END
END A6
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER ME4 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER ME3 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER ME2 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER ME1 ;
  RECT 267.900 0.000 269.020 1.120 ;
 END
END A5
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER ME4 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER ME3 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER ME2 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER ME1 ;
  RECT 262.320 0.000 263.440 1.120 ;
 END
END A4
PIN A9
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 249.300 0.000 250.420 1.120 ;
  LAYER ME4 ;
  RECT 249.300 0.000 250.420 1.120 ;
  LAYER ME3 ;
  RECT 249.300 0.000 250.420 1.120 ;
  LAYER ME2 ;
  RECT 249.300 0.000 250.420 1.120 ;
  LAYER ME1 ;
  RECT 249.300 0.000 250.420 1.120 ;
 END
END A9
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 243.720 0.000 244.840 1.120 ;
  LAYER ME4 ;
  RECT 243.720 0.000 244.840 1.120 ;
  LAYER ME3 ;
  RECT 243.720 0.000 244.840 1.120 ;
  LAYER ME2 ;
  RECT 243.720 0.000 244.840 1.120 ;
  LAYER ME1 ;
  RECT 243.720 0.000 244.840 1.120 ;
 END
END A8
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME4 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME3 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME2 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME1 ;
  RECT 237.520 0.000 238.640 1.120 ;
 END
END A7
PIN DIA3
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 161.260 0.000 162.380 1.120 ;
  LAYER ME4 ;
  RECT 161.260 0.000 162.380 1.120 ;
  LAYER ME3 ;
  RECT 161.260 0.000 162.380 1.120 ;
  LAYER ME2 ;
  RECT 161.260 0.000 162.380 1.120 ;
  LAYER ME1 ;
  RECT 161.260 0.000 162.380 1.120 ;
 END
END DIA3
PIN DOA3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 147.620 0.000 148.740 1.120 ;
  LAYER ME4 ;
  RECT 147.620 0.000 148.740 1.120 ;
  LAYER ME3 ;
  RECT 147.620 0.000 148.740 1.120 ;
  LAYER ME2 ;
  RECT 147.620 0.000 148.740 1.120 ;
  LAYER ME1 ;
  RECT 147.620 0.000 148.740 1.120 ;
 END
END DOA3
PIN DIA2
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER ME4 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER ME3 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER ME2 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER ME1 ;
  RECT 133.980 0.000 135.100 1.120 ;
 END
END DIA2
PIN DOA2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 120.960 0.000 122.080 1.120 ;
  LAYER ME4 ;
  RECT 120.960 0.000 122.080 1.120 ;
  LAYER ME3 ;
  RECT 120.960 0.000 122.080 1.120 ;
  LAYER ME2 ;
  RECT 120.960 0.000 122.080 1.120 ;
  LAYER ME1 ;
  RECT 120.960 0.000 122.080 1.120 ;
 END
END DOA2
PIN DIA1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER ME4 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER ME3 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER ME2 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER ME1 ;
  RECT 52.760 0.000 53.880 1.120 ;
 END
END DIA1
PIN DOA1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER ME4 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER ME3 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER ME2 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER ME1 ;
  RECT 39.740 0.000 40.860 1.120 ;
 END
END DOA1
PIN DIA0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER ME4 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER ME3 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER ME2 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER ME1 ;
  RECT 26.100 0.000 27.220 1.120 ;
 END
END DIA0
PIN DOA0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER ME4 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER ME3 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER ME2 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER ME1 ;
  RECT 12.460 0.000 13.580 1.120 ;
 END
END DOA0
OBS
  LAYER ME1 SPACING 0.280 ;
  RECT 0.000 0.140 544.980 349.860 ;
  LAYER ME2 SPACING 0.320 ;
  RECT 0.000 0.140 544.980 349.860 ;
  LAYER ME3 SPACING 0.320 ;
  RECT 0.000 0.140 544.980 349.860 ;
  LAYER ME4 SPACING 0.600 ;
  RECT 0.000 0.140 544.980 349.860 ;
  LAYER VI1 ;
  RECT 0.000 0.140 544.980 349.860 ;
  LAYER VI2 ;
  RECT 0.000 0.140 544.980 349.860 ;
  LAYER VI3 ;
  RECT 0.000 0.140 544.980 349.860 ;
END
END W1024_B8_BM2
END LIBRARY



