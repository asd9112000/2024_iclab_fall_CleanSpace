../00_TESTBED/TA_PATTERN.sv